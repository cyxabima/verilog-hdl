module ground(output zero);
    assign zero = 0;
endmodule