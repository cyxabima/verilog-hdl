module and_gate(output y,input a,b);
    assign y = a & b; //  & bit wise or && logical or since we have only one bit so both are same
endmodule