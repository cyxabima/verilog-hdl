module vcc(output one);
    assign one = 1;
endmodule